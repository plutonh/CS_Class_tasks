`timescale 1ns / 1ps

module assignment_1(
	input [31:0] a, b,
	output [31:0] c, d
	);
	
	assign c = a;
	assign d = b;
endmodule