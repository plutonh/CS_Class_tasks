`timescale 1ns / 1ps

module Branch_Prediction(
    );


endmodule
